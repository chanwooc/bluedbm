// Copyright (c) 2013 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import CtrlMux::*;
import Portal::*;
import Leds::*;
import ConnectalMemory::*;
import MemTypes::*;
import MemServer::*;
import MMU::*;

import HostInterface::*;

// generated by tool
import FlashRequest::*;
import FlashIndication::*;

// generated by tool: hopefully only this part will change
import MemServerRequest::*;
import MMURequest::*;
import MemServerIndication::*;
import MMUIndication::*;

`ifndef BSIM
import Xilinx       :: *;
import XilinxCells ::*;
import DefaultValue    :: *;
`endif
import Clocks :: *;


// defined by user
import Main::*;

import AuroraCommon::*;

typedef enum {FlashIndicationH2S, FlashRequestS2H, HostMemServerIndicationH2S, HostMemServerRequestS2H, HostMMURequestS2H, HostMMUIndicationH2S
	} IfcNames deriving (Eq,Bits);

interface Top_Pins;
	interface Aurora_Pins#(4) aurora_fmc1;
	interface Aurora_Clock_Pins aurora_clk_fmc1;
endinterface

//typedef 128 DataBusWidth;

module mkConnectalTop#(Clock clk250, Reset rst250) (ConnectalTop#(PhysAddrWidth,DataBusWidth,Top_Pins,NumberOfMasters))
   provisos (Add#(0,128,DataBusWidth),Add#(1,0,NumberOfMasters));

	
	Clock curClk <- exposeCurrentClock;
	Reset curRst <- exposeCurrentReset;

	/////////////////////////////////////////

   FlashIndicationProxy flashIndicationProxy <- mkFlashIndicationProxy(FlashIndicationH2S);

   MainIfc hwmain <- mkMain(flashIndicationProxy.ifc, clk250, rst250);
   FlashRequestWrapper flashRequestWrapper <- mkFlashRequestWrapper(FlashRequestS2H,hwmain.request);

   //Vector#(1,  MemReadClient#(DataBusWidth))   readClients = cons(hwmain.dmaReadClient, nil);
   //Vector#(1, MemWriteClient#(DataBusWidth))  writeClients = cons(hwmain.dmaWriteClient, nil);
   
   let readClients = hwmain.dmaReadClient;
   let writeClients = hwmain.dmaWriteClient;

   
   MMUIndicationProxy hostMMUIndicationProxy <- mkMMUIndicationProxy(HostMMUIndicationH2S);
   MMU#(PhysAddrWidth) hostMMU <- mkMMU(0, True, hostMMUIndicationProxy.ifc);
   MMURequestWrapper hostMMURequestWrapper <- mkMMURequestWrapper(HostMMURequestS2H, hostMMU.request);

   MemServerIndicationProxy hostMemServerIndicationProxy <- mkMemServerIndicationProxy(HostMemServerIndicationH2S);
   MemServer#(PhysAddrWidth,DataBusWidth,1) dma <- mkMemServer(readClients, writeClients, cons(hostMMU,nil), hostMemServerIndicationProxy.ifc);
   MemServerRequestWrapper hostMemServerRequestWrapper <- mkMemServerRequestWrapper(HostMemServerRequestS2H, dma.request);

   Vector#(6,StdPortal) portals;
   portals[0] = flashRequestWrapper.portalIfc;
   portals[1] = flashIndicationProxy.portalIfc; 
   portals[2] = hostMemServerRequestWrapper.portalIfc;
   portals[3] = hostMemServerIndicationProxy.portalIfc; 
   portals[4] = hostMMURequestWrapper.portalIfc;
   portals[5] = hostMMUIndicationProxy.portalIfc;
   
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;

	interface Top_Pins pins;
		interface Aurora_Pins aurora_fmc1 = hwmain.aurora_fmc1;
		interface Aurora_Clock_Pins aurora_clk_fmc1 = hwmain.aurora_clk_fmc1;
	endinterface
endmodule


