
typedef enum {FlashIndicationH2S, FlashRequestS2H, PlatformIfcNames_MemServerIndicationH2S, PlatformIfcNames_MemServerRequestS2H, PlatformIfcNames_MMURequestS2H, PlatformIfcNames_MMUIndicationH2S
	} IfcNames deriving (Eq,Bits);

